version https://git-lfs.github.com/spec/v1
oid sha256:a451df9f967cc624ba952d79ecb37f9ed0fb05437f4a5b2d169d2959381e68df
size 63005

version https://git-lfs.github.com/spec/v1
oid sha256:a0faf8ef7d33c4f794633bbaac16a747b69f7c9eb88e0871d9b56041fdcc195f
size 131533

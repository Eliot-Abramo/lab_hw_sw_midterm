version https://git-lfs.github.com/spec/v1
oid sha256:45664b6ad2f92ef23692c5d071b932cf85260c94e24b028363a37e45b48da88e
size 1500

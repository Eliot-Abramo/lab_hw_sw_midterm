version https://git-lfs.github.com/spec/v1
oid sha256:b8b6bece785281b3ce3ca2a351b5bee17b97b0cdc2cc4bf8bcd8a3c24e240343
size 1498

version https://git-lfs.github.com/spec/v1
oid sha256:a26922b433a3acd83c13c9e27e9a63d51db8895d755fb2f14010250ad8e9be29
size 22922

version https://git-lfs.github.com/spec/v1
oid sha256:00e3cdd0468258958cc1802a6dc4ef662a2659e29cf91358d409f203c75df8fd
size 94742

version https://git-lfs.github.com/spec/v1
oid sha256:b51e8b914b45510d6c7a369bf181f6fc2db18cbffbe49c2e40366cb920e0e609
size 1480

version https://git-lfs.github.com/spec/v1
oid sha256:0acab6e3ffc785102f79fe18f242746afec5b606941a1f41919f2bf09129b901
size 40102

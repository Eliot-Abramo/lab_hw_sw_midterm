version https://git-lfs.github.com/spec/v1
oid sha256:03d0fdc03a340ce3bfca9c7e58741efb4e00872f143099306c1c46b17fcfd5dc
size 1500

version https://git-lfs.github.com/spec/v1
oid sha256:f795b3e2115489a59437713ee6a198c008e5fe88d910c07610d3f63176293534
size 1964

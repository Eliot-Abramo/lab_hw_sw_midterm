version https://git-lfs.github.com/spec/v1
oid sha256:b0e7d6bc2b5fb81a8fbc8961a80d8c9880f81c230b7cd8a07ce0f544b57745c6
size 2311

version https://git-lfs.github.com/spec/v1
oid sha256:8bb4d5ce949e7f5d6b2dc1647a45f14c98dc906ae057146414370560762d1b15
size 1964

version https://git-lfs.github.com/spec/v1
oid sha256:785bc24cdc43249ad6d7750255397740c50ed0a570b55b8d21e31f48228ed212
size 1061

version https://git-lfs.github.com/spec/v1
oid sha256:305d9523112079e732cea175386a63ca99c3f563acc20fa6f341198ea5190fbf
size 2074

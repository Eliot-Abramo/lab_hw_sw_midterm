version https://git-lfs.github.com/spec/v1
oid sha256:0fc60a2b6437cc5155d38dc3c996d3aa12058ac394093aa24b75b0971259094c
size 1610

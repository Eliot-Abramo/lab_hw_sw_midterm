version https://git-lfs.github.com/spec/v1
oid sha256:ca7024d01faff9ff9cde1ea916f4638fc4a777053ca2b6123534469c15d5dd38
size 26937

version https://git-lfs.github.com/spec/v1
oid sha256:a36d4f73331672601480c00b173e70d347629392e28b260982df6029e60a0093
size 45023

version https://git-lfs.github.com/spec/v1
oid sha256:7691f41bc8f6e5810a754106ea447c86457827e468c39ae6b40044696835e1f5
size 146813

version https://git-lfs.github.com/spec/v1
oid sha256:3625ef933e98bd3912f91b3023b84b66f689c9e9ca9151929601462629a669ed
size 43049

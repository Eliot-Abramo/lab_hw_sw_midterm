version https://git-lfs.github.com/spec/v1
oid sha256:8932cfb8246ed9567270184578d69f788db6e7e07744545cf4f5eaadd56a03df
size 1081

version https://git-lfs.github.com/spec/v1
oid sha256:7863d3faa773ec30da3f7e6995782615d350da60c12f33e667b8fe6f90883d24
size 2321

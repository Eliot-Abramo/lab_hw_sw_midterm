version https://git-lfs.github.com/spec/v1
oid sha256:c531c9d28687c9fe8716ee451a629b872510ae209b17a1d3c4355705705ae34c
size 2342

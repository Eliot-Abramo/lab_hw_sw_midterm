version https://git-lfs.github.com/spec/v1
oid sha256:7d854f30d6fee043e53024d9ad05e0c3824b8bb60604d5bfb5bdfd6a9a03496e
size 38399

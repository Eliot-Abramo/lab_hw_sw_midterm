version https://git-lfs.github.com/spec/v1
oid sha256:8762aac641d9e69b8e8233f90ec89b00a169f6efd03eaaa84e04409f5db9d068
size 1776

version https://git-lfs.github.com/spec/v1
oid sha256:32b0fb9d7ef5f8ce733059edf212d1a0e2b2fc1beca3cc65225164d83579ba43
size 56878

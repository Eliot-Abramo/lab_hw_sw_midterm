version https://git-lfs.github.com/spec/v1
oid sha256:97929fb0ba870bb000fae49224861e5ecc2961a6d37ae7adf9c7d16cf34fa216
size 146813

version https://git-lfs.github.com/spec/v1
oid sha256:ca78751e22e75534ef154d026af1cb1d2c4b6d50d912a91caa0629be1b5ecf07
size 1081

version https://git-lfs.github.com/spec/v1
oid sha256:8fa61e8d31ff0ce5bf51166d4ffd4c9409e02b29dc91f53c2fff5b94fcb04138
size 2082

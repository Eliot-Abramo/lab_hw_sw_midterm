version https://git-lfs.github.com/spec/v1
oid sha256:9c98f429d7b048e6dc7f945f8efd8505c1c62f87d8d465167d7647ed8692d708
size 146728

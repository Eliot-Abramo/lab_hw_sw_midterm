version https://git-lfs.github.com/spec/v1
oid sha256:cb504daddaa771f55f20a82938dc07f37542aa6ddd40693aac95aa75111dcb73
size 94472

version https://git-lfs.github.com/spec/v1
oid sha256:462d15e175834fe2cf05b3d2f322a399416ce2dbaa75d9ac5a2bba9538774cdd
size 45010

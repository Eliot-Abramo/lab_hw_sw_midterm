version https://git-lfs.github.com/spec/v1
oid sha256:fa1de3962e47000d73b3061642f0313613c2b8ac2518a3d0109e014af2ee0dc6
size 1500

version https://git-lfs.github.com/spec/v1
oid sha256:613cf9effe62b09c9a03f009dad66f8ffe0f55de7fde30cf406090b15774918f
size 3014

version https://git-lfs.github.com/spec/v1
oid sha256:1eec30555ad3d0089f7d84701d8438a803e3bc421523a18c8b9184d114f9f3b4
size 119955

version https://git-lfs.github.com/spec/v1
oid sha256:546e96c7ee0a1b30099d48d28d1a0ff82a1ddf5a3c925d8ca77b0ecb2629480e
size 80260

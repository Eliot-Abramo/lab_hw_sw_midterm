version https://git-lfs.github.com/spec/v1
oid sha256:1fc996c7e4b697ee26b928442422909d6940feb6e1a6c36eebc8ad41202279ac
size 56902

version https://git-lfs.github.com/spec/v1
oid sha256:85b6e4076717cb9df137bdf1ee90d7e88567d4ba8c0c32eb54f9bcd7c7081aee
size 40418

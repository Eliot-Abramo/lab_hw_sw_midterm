version https://git-lfs.github.com/spec/v1
oid sha256:39b0319120899e1f8e712aa6d6bb54f403302ddfa131c8934cb7aaff2fafb699
size 1944

version https://git-lfs.github.com/spec/v1
oid sha256:b9eceec78d3102e5f48316918d6ead2ae00a70d76fce227272efd465ab5ab68e
size 2315

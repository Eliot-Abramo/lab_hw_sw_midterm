version https://git-lfs.github.com/spec/v1
oid sha256:b0899ebd33ca8e40f5ed736ef0ca2e093013589e9474c613e08db852e63bb521
size 1087

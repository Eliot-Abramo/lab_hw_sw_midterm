version https://git-lfs.github.com/spec/v1
oid sha256:04086430c8ce78eca3ba206bdf5ff1b933b852b4165befeaf7ef909f7a7269bf
size 43103

version https://git-lfs.github.com/spec/v1
oid sha256:0b3a7af146ce74dd3243868b30f032a962168e670ceac9f568bad2dad334d55d
size 2070

version https://git-lfs.github.com/spec/v1
oid sha256:d51f2afce710779320d484024137f87021b01a9af198c4236548890d4718b167
size 99647

version https://git-lfs.github.com/spec/v1
oid sha256:d0697da4ca84a69f081f4c2104b674b72ed1ac9a9d9973a070fe675913d9ca9f
size 193991

version https://git-lfs.github.com/spec/v1
oid sha256:f6047af2ec0c81ae92f32596747f5ceac686de7f3672adea8e8b3fe2ed2547e2
size 25312

version https://git-lfs.github.com/spec/v1
oid sha256:09b3aa54f8639e9d7f69444fcf858486f3840dad6b19093fcc40730183b79470
size 12126

version https://git-lfs.github.com/spec/v1
oid sha256:ab983198ced4240f1ee30faaebabe1b87f1b3174db8b9b01fc1a5fabb17a36be
size 56937

version https://git-lfs.github.com/spec/v1
oid sha256:c9df6703e983129726170ee3000a10692853a7ecef8ef2b39de30496fb3a2478
size 40365

version https://git-lfs.github.com/spec/v1
oid sha256:95edea9f38315471f7ececb77bc7eb4b15be4f27c3f71f4e3923bc05ba0469d8
size 164698

version https://git-lfs.github.com/spec/v1
oid sha256:433a99561b658dafc8d7925fa81cada4d190729eeb070f61a87a25732e1940d6
size 3265

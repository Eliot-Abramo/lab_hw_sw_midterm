version https://git-lfs.github.com/spec/v1
oid sha256:e1d9fc167d63f233baef5e1821ac9e665d49db426b066d17aadc8a004e7a1106
size 146813

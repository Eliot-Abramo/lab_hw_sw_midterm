version https://git-lfs.github.com/spec/v1
oid sha256:0020d01ba7361d3bbeb35b620348395224aa12b869419effb639e91f4b48fa4c
size 55661

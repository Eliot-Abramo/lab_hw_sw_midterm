version https://git-lfs.github.com/spec/v1
oid sha256:b2120e03792c9aaaa33ce0d1902cc583c18e42edc62806960e5747ee279c64dd
size 146813

version https://git-lfs.github.com/spec/v1
oid sha256:fd3c0c901580b9faf0978a90c31302c0715c82ddfec0b3d8aa750cc293777d36
size 45007

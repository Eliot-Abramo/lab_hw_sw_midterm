version https://git-lfs.github.com/spec/v1
oid sha256:5195bdbc465e400ad157ee9e73b9379e60ef4c0895716e29d55fbd6a2e58e5d4
size 42867

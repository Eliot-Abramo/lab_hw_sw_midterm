version https://git-lfs.github.com/spec/v1
oid sha256:400b0533f0d255c2e009a6a0cbbaf1d9117a478c54489e65b19329fde9222070
size 1500

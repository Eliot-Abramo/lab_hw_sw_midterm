version https://git-lfs.github.com/spec/v1
oid sha256:8b0b396774e7c99ce7b5bc974e552340a1093a9de6a681033813b5edb58bb8dd
size 44245

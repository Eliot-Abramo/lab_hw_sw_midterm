version https://git-lfs.github.com/spec/v1
oid sha256:a6e934a7f04c33a4903632ea885b0c4aeee6a116a5cefb5981e71533e40cac44
size 2327

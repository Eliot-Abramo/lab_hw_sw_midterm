version https://git-lfs.github.com/spec/v1
oid sha256:4fd5adaaa6190698bc08734e19eb5b8ebd19d6f65a59bd240db7fe0b1d15c07f
size 133486

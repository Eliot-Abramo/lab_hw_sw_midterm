version https://git-lfs.github.com/spec/v1
oid sha256:07167dcb0db4b7cb8b9dee66a6d6cfb50e2af93179f9afcfa7824b6aa4be1948
size 101834

version https://git-lfs.github.com/spec/v1
oid sha256:1f5e803a6a008d0630b15b942f559924597b9424089d3678b54ab503212b696e
size 103759

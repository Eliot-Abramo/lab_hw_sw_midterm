version https://git-lfs.github.com/spec/v1
oid sha256:df698c387562a75f8955689f8f9036fcbcf7047e869eda7b1c40500e268bdb1c
size 1964

version https://git-lfs.github.com/spec/v1
oid sha256:0130bc02e50640a19a2fa1a5b3252c2fd2897c0b1225338fd3e868c735a9fb72
size 276477
